--addi rd, rs1, imm
imm[12bits] rs1 000 rd 0010011                    ---- 010000000000 00010 000 00010 0010011
--sw
imm[11:5] rs2 rs1 010 imm[4:0] 0100011
--jal x0, label
imm[20|10:1|11|19:12] rd 1101111
--slli
imm(12bits) rs1 001 rd 0010011
---add
0000000 rs2 rs1 000 rd 0110011
--bge
imm[12|10:5] rs2 rs1 101 imm[4:1|11] 1100011
--lw
imm(12bits) rs1 010 rd 0000011
--sub
0100000 rs2 rs1 000 rd 0110011
--blt
imm[12|10:5] rs2 rs1 100 imm[4:1|11] 1100011
--jalr x0, 0(x1)
imm(12bits) rs1 000 rd 1100111
-------------------------------------------------------------------------------
01000000000000010000000100010011     -- sp to 1024
01000000000001000000010000010011     -- s0 to 1024


111111010000 00010 000 00010 0010011  -- addi	sp,sp,-48
0000001 01000 00010 010 01100 0100011      --sw	s0,44(sp)
000000110000 00010 000 01000 0010011      --addi	s0,sp,48
000000000011 01111 000 01111 0010011     -- li	a5,3         addi a5,a5,3

00000000001101111000011110010011
  0100011110001101

1111110 01111 01000 010 10000 0100011      -- sw	a5,-48(s0)
000000000101 01111 000 01111 0010011     -- 	li	a5,5
1111110 01111 01000 010 10100 0100011      -- sw	a5,-44(s0)
000000000001 01111 000 01111 0010011    -- li	a5,1
1111110 01111 01000 010 11000 0100011      -- sw	a5,-40(s0)
000000000010 01111 000 01111 0010011    -- li	a5,2
1111110 01111 01000 010 11100 0100011      -- sw	a5,-36(s0)
000000000100 01111 000 01111 0010011    -- li	a5,4
1111111 01111 01000 010 00000 0100011      -- sw	a5,-32(s0)
1111111 00000 01000 010 01100 0100011    -- 	sw	zero,-20(s0)
00000110010000000000 00000 1101111  -- 	j	.L2    --jal x0, 200  (immediate encoded here is 000000000000001100100 It is 100-decimal bec it gets shifted by <<1 in the datapath)
1111111 00000 01000 010 01000 0100011    -- 	sw	zero,-24(s0)                             
00000101000000000000 00000 1101111  -- 	j	.L3    --jal x0, 160
111111101000 01000 010 01111 0000011 -- lw a5,-24(s0)
000000000010 01111 001 01111 0010011  --	slli	a5,a5,2
111111110000 01000 000 01110 0010011  -- 	addi	a4,s0,-16
0000000 01111 01110 000 01111 0110011 -- 	add	a5,a4,a5
111111100000 01111 010 01110 0000011 -- lw a4,-32(a5)
111111101000 01000 010 01111 0000011 -- lw a5,-24(s0)
000000000001 01111 000 01111 0010011  -- 	addi	a5,a5,1
000000000010 01111 001 01111 0010011  --	slli	a5,a5,2
111111110000 01000 000 01101 0010011  -- 	addi	a3,s0,-16
0000000 01111 01101 000 01111 0110011 -- 	add	a5,a3,a5
111111100000 01111 010 01111 0000011 -- 	lw	a5,-32(a5)
0000001 01110 01111 101 10010 1100011  -- bge	a5,a4,.L4

--#load arr[j] a5
lw	a5,-24(s0)
slli	a5,a5,2
addi	a4,s0,-16
add	a5,a4,a5
lw	a5,-32(a5)








	


